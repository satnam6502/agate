module adder8(
  input  logic cin,
  input  logic [7:0] x,
  input  logic [7:0] y,
  output logic [7:0] sum,
  output logic cout);
  logic net40;
  logic net39;
  logic net38;
  logic net37;
  logic net36;
  logic net35;
  logic net34;
  logic net33;
  logic net32;
  logic net31;
  logic net30;
  logic net29;
  logic net28;
  logic net27;
  logic net26;
  logic net25;
  logic net24;
  logic net23;
  logic net22;
  logic net21;
  logic net20;
  logic net19;
  logic net18;
  logic net17;
  logic net16;
  logic net15;
  logic net14;
  logic net13;
  logic net12;
  logic net11;
  logic net10;
  logic net9;
  logic net8;
  logic net7;
  logic net6;
  logic net5;
  logic net4;
  logic net3;
  logic net2;
  logic net1;
  logic net0;

  logic [7:0] vec0;
  logic [7:0] vec1;
  assign cout = net40;
  assign sum = '{net38, net33, net28, net23, net18, net13, net8, net3};
  or (net40, net37, net39);
  and (net39, net36, net35);
  xor (net38, net36, net35);
  and (net37, vec0[7], vec1[7]);
  xor (net36, vec0[7], vec1[7]);
  or (net35, net32, net34);
  and (net34, net31, net30);
  xor (net33, net31, net30);
  and (net32, vec0[6], vec1[6]);
  xor (net31, vec0[6], vec1[6]);
  or (net30, net27, net29);
  and (net29, net26, net25);
  xor (net28, net26, net25);
  and (net27, vec0[5], vec1[5]);
  xor (net26, vec0[5], vec1[5]);
  or (net25, net22, net24);
  and (net24, net21, net20);
  xor (net23, net21, net20);
  and (net22, vec0[4], vec1[4]);
  xor (net21, vec0[4], vec1[4]);
  or (net20, net17, net19);
  and (net19, net16, net15);
  xor (net18, net16, net15);
  and (net17, vec0[3], vec1[3]);
  xor (net16, vec0[3], vec1[3]);
  or (net15, net12, net14);
  and (net14, net11, net10);
  xor (net13, net11, net10);
  and (net12, vec0[2], vec1[2]);
  xor (net11, vec0[2], vec1[2]);
  or (net10, net7, net9);
  and (net9, net6, net5);
  xor (net8, net6, net5);
  and (net7, vec0[1], vec1[1]);
  xor (net6, vec0[1], vec1[1]);
  or (net5, net2, net4);
  and (net4, net1, net0);
  xor (net3, net1, net0);
  and (net2, vec0[0], vec1[0]);
  xor (net1, vec0[0], vec1[0]);
  assign vec1 = y;
  assign vec0 = x;
  assign net0 = cin;
endmodule: adder8